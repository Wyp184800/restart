module	flash_top